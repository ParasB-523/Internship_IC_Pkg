VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO C4BUMP
	CLASS COVER BUMP ;
	ORIGIN 0 0 ;
	SIZE 70 BY 70 ;
	SYMMETRY X Y ;
	PIN PAD
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER metal1 ;
		    		POLYGON 20.5025 0 49.4975 0 70 20.5025 70 49.4975 49.4975 70 20.5025 70 0 49.4975 0 20.5025 ;
		  	LAYER via1 ;
		    		RECT 25 23 45 47 ;
		  	LAYER metal2 ;
		    		RECT 22 20 48 50 ;
		END
	END PAD
	OBS
	  	LAYER metal2 SPACING 0.000 ;
	    		RECT 20 18 50 19 ;
	    		RECT 20 51 50 52 ;
	    		RECT 20 18 21 51 ;
	    		RECT 49 18 50 51 ;
	END
END C4BUMP

END LIBRARY