VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO UBUMP
	CLASS COVER BUMP ;
	ORIGIN 0 0 ;
	SIZE 22.5 BY 22.5 ;
	SYMMETRY X Y ;
	PIN PAD
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER metal6 ;
				POLYGON 6.59 0 15.91 0 22.5 6.59 22.5 15.91 15.91 22.5 6.59 22.5 0 15.91 0 6.59 ; 
		END
	END PAD
	OBS
		LAYER via5 SPACING 0.000 ;
			POLYGON 6.59 2 15.91 2 20.5 6.59 20.5 15.91 15.91 20.5 6.59 20.5 2 15.91 2 6.59 ; 
	END
END UBUMP

END LIBRARY